module unmasked_aes_sbox(in, out);
  input [7:0] in;
  output [7:0] out;
  wire [7:0] in;
  wire [7:0] out;
  wire n_4, n_7, n_8, n_9, n_11, n_13, n_15, n_16;
  wire n_19, n_20, n_21, n_23, n_24, n_25, n_27, n_28;
  wire n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52;
  wire n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60;
  wire n_61, n_62, n_63, n_64, n_65, n_66, n_67, n_68;
  wire n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84;
  wire n_85, n_86, n_87, n_88, n_89, n_90, n_91, n_92;
  wire n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100;
  wire n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108;
  wire n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
  wire n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124;
  wire n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132;
  wire n_133, n_134, n_135, n_136, n_137, n_138, n_139, n_140;
  wire n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148;
  wire n_149, n_150, n_151, n_152, n_153, n_154, n_155, n_156;
  wire n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164;
  wire n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172;
  wire n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180;
  wire n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188;
  wire n_189, n_190, n_192, n_193, n_195, n_196, n_197, n_198;
  wire n_199, n_200, n_201;
  xnor XNOR2_g2018(out[7], n_181, out[5]);
  xnor XNOR2_g2019(out[4], n_178, n_200);
  xnor XNOR2_g2020(out[2], n_198, n_190);
  xnor XNOR2_g2022(out[1], n_195, n_201);
  xnor XNOR2_g2021(out[0], n_192, n_199);
  xnor XNOR2_g2023(out[5], n_196, n_201);
  xnor XNOR2_g2026(n_200, n_197, n_199);
  xnor XNOR2_g2027(n_198, n_180, n_197);
  xnor XNOR2_g2025(n_196, n_188, n_193);
  xnor XNOR2_g2024(n_195, n_193, out[3]);
  xnor XNOR2_g2028(n_192, n_189, out[3]);
  xnor XNOR2_g2034(n_197, n_187, n_173);
  xnor XNOR2_g2032(out[6], n_186, n_201);
  xnor XNOR2_g2030(n_193, n_179, n_190);
  xnor XNOR2_g2033(n_189, n_174, n_183);
  xnor XNOR2_g2031(n_199, n_185, n_175);
  xnor XNOR2_g2029(n_188, n_177, n_172);
  not NOT1_g2035(n_187, n_186);
  xnor XNOR2_g2041(n_185, n_117, n_184);
  xnor XNOR2_g2037(n_186, n_139, n_182);
  xnor XNOR2_g2039(n_201, n_127, n_184);
  xnor XNOR2_g2042(n_183, n_168, n_182);
  xnor XNOR2_g2043(n_181, n_151, n_180);
  xnor XNOR2_g2036(n_179, n_161, n_178);
  xnor XNOR2_g2038(out[3], n_160, n_176);
  xnor XNOR2_g2040(n_177, n_176, n_190);
  xnor XNOR2_g2049(n_182, n_145, n_166);
  xnor XNOR2_g2050(n_178, n_116, n_171);
  xnor XNOR2_g2045(n_175, n_174, n_167);
  xnor XNOR2_g2048(n_184, n_165, n_169);
  xnor XNOR2_g2046(n_180, n_164, n_170);
  xnor XNOR2_g2044(n_173, n_162, n_172);
  xnor XNOR2_g2047(n_176, n_158, n_163);
  xnor XNOR2_g2051(n_171, n_118, n_148);
  xnor XNOR2_g2052(n_170, n_126, n_153);
  xnor XNOR2_g2053(n_169, n_150, n_141);
  xnor XNOR2_g2054(n_168, n_142, n_159);
  xnor XNOR2_g2055(n_167, n_156, n_144);
  xnor XNOR2_g2057(n_166, n_157, n_123);
  xnor XNOR2_g2058(n_165, n_135, n_114);
  xnor XNOR2_g2059(n_164, n_113, n_132);
  xnor XNOR2_g2056(n_172, n_120, n_124);
  xnor XNOR2_g2061(n_163, n_130, n_146);
  xnor XNOR2_g2060(n_162, n_160, n_161);
  xnor XNOR2_g2062(n_174, n_137, n_121);
  xnor XNOR2_g2063(n_190, n_129, n_125);
  nand NAND2_g2086(n_159, n_147, n_155);
  nand NAND2_g2083(n_158, n_149, n_152);
  nand NAND2_g2081(n_157, n_154, n_44);
  nand NAND2_g2091(n_156, n_154, n_155);
  nand NAND2_g2065(n_153, n_154, n_152);
  not NOT1_g2064(n_151, n_161);
  nand NAND2_g2092(n_150, n_149, n_155);
  nand NAND2_g2072(n_148, n_147, n_152);
  nor NOR2_g2084(n_146, n_131, n_140);
  nor NOR2_g2085(n_145, n_143, n_136);
  nor NOR2_g2087(n_144, n_143, n_134);
  nand NAND2_g2088(n_142, n_138, n_35);
  nor NOR2_g2089(n_141, n_143, n_140);
  nand NAND2_g2090(n_139, n_138, n_155);
  nor NOR2_g2093(n_137, n_133, n_136);
  nor NOR2_g2094(n_135, n_133, n_134);
  nor NOR2_g2096(n_132, n_131, n_134);
  nor NOR2_g2066(n_130, n_128, n_134);
  nor NOR2_g2068(n_129, n_128, n_140);
  nor NOR2_g2069(n_127, n_122, n_136);
  nor NOR2_g2070(n_126, n_119, n_136);
  nor NOR2_g2071(n_125, n_131, n_136);
  nand NAND2_g2073(n_124, n_138, n_152);
  nor NOR2_g2074(n_123, n_122, n_134);
  nor NOR2_g2075(n_121, n_122, n_140);
  nor NOR2_g2077(n_120, n_119, n_134);
  nor NOR2_g2078(n_118, n_119, n_140);
  nor NOR2_g2080(n_161, n_128, n_136);
  nor NOR2_g2095(n_117, n_133, n_115);
  nor NOR2_g2082(n_116, n_131, n_115);
  not NOT1_g2097(n_149, n_136);
  not NOT1_g2098(n_147, n_134);
  nor NOR2_g2076(n_114, n_122, n_115);
  nor NOR2_g2067(n_113, n_128, n_115);
  nor NOR2_g2079(n_160, n_119, n_115);
  not NOT1_g2102(n_154, n_140);
  nor NOR2_g2099(n_136, n_77, n_111);
  nor NOR2_g2100(n_134, n_112, n_109);
  not NOT1_g2101(n_138, n_115);
  nor NOR2_g2104(n_140, n_106, n_110);
  nor NOR2_g2103(n_115, n_112, n_108);
  nand NAND2_g2105(n_111, n_105, n_104);
  nand NAND2_g2107(n_110, n_103, n_84);
  nand NAND2_g2108(n_109, n_107, n_102);
  nand NAND2_g2106(n_108, n_101, n_76);
  nor NOR2_g2111(n_107, n_94, n_80);
  nor NOR2_g2112(n_106, n_96, n_95);
  nor NOR2_g2113(n_105, n_98, n_86);
  nor NOR2_g2114(n_104, n_100, n_88);
  nand NAND2_g2115(n_103, n_99, n_93);
  nor NOR2_g2109(n_102, n_92, n_89);
  nor NOR2_g2110(n_101, n_82, n_90);
  nor NOR2_g2117(n_100, n_81, n_75);
  nand NAND2_g2126(n_99, n_91, n_97);
  nor NOR2_g2127(n_98, n_96, n_97);
  nand NAND2_g2130(n_95, n_71, n_87);
  nor NOR2_g2119(n_94, n_93, n_97);
  nor NOR2_g2120(n_92, n_96, n_91);
  nor NOR2_g2118(n_90, n_91, n_85);
  not NOT1_g2116(n_89, n_79);
  nor NOR2_g2121(n_88, n_87, n_91);
  nor NOR2_g2129(n_86, n_83, n_85);
  nand NAND2_g2125(n_84, n_70, n_83);
  not NOT1_g2124(n_82, n_73);
  nor NOR2_g2132(n_112, n_81, n_69);
  nor NOR2_g2122(n_80, n_78, n_85);
  nand NAND2_g2123(n_79, n_77, n_78);
  nand NAND2_g2128(n_76, n_85, n_74);
  nand NAND2_g2133(n_75, n_72, n_74);
  nand NAND2_g2131(n_73, n_77, n_72);
  not NOT1_g2136(n_71, n_83);
  nand NAND2_g2134(n_97, n_68, n_74);
  not NOT1_g2137(n_70, n_85);
  nand NAND2_g2135(n_91, n_72, n_78);
  nand NAND2_g2138(n_69, n_93, n_68);
  nand NAND2_g2140(n_83, n_68, n_78);
  nor NOR2_g2139(n_77, n_87, n_96);
  not NOT1_g2142(n_74, n_78);
  nand NAND2_g2141(n_85, n_96, n_87);
  not NOT1_g2143(n_81, n_96);
  xnor XNOR2_g2144(n_78, n_67, n_48);
  not NOT1_g2146(n_68, n_72);
  not NOT1_g2147(n_93, n_87);
  xnor XNOR2_g2145(n_96, n_65, n_62);
  xnor XNOR2_g2148(n_72, n_66, n_60);
  xnor XNOR2_g2149(n_87, n_64, n_58);
  xnor XNOR2_g2151(n_67, n_49, n_59);
  xnor XNOR2_g2150(n_66, n_39, n_61);
  xnor XNOR2_g2152(n_65, n_57, n_63);
  xnor XNOR2_g2153(n_64, n_11, n_63);
  xnor XNOR2_g2154(n_62, n_19, n_61);
  xnor XNOR2_g2155(n_60, n_56, n_47);
  xnor XNOR2_g2159(n_59, n_29, n_55);
  xnor XNOR2_g2156(n_58, n_51, n_37);
  xnor XNOR2_g2157(n_63, n_28, n_54);
  xnor XNOR2_g2158(n_57, n_36, n_52);
  xnor XNOR2_g2160(n_61, n_7, n_53);
  xnor XNOR2_g2167(n_56, n_46, n_34);
  nor NOR2_g2162(n_55, n_42, n_50);
  xnor XNOR2_g2166(n_54, n_41, n_24);
  xnor XNOR2_g2168(n_53, n_43, n_30);
  nand NAND2_g2161(n_52, n_155, n_38);
  nand NAND2_g2163(n_51, n_155, n_45);
  not NOT1_g2169(n_50, n_155);
  xnor XNOR2_g2164(n_49, in[3], n_27);
  xnor XNOR2_g2165(n_48, n_31, n_47);
  nand NAND2_g2178(n_46, n_44, n_45);
  nand NAND2_g2170(n_155, n_40, n_33);
  nor NOR2_g2176(n_43, n_42, n_133);
  nor NOR2_g2183(n_41, n_32, n_133);
  not NOT1_g2173(n_40, n_39);
  xnor XNOR2_g2171(n_152, n_143, n_38);
  xnor XNOR2_g2172(n_131, n_143, n_37);
  nand NAND2_g2180(n_36, n_35, n_45);
  nand NAND2_g2184(n_34, n_35, n_38);
  not NOT1_g2186(n_44, n_133);
  nand NAND2_g2174(n_33, n_32, in[4]);
  nor NOR2_g2182(n_31, n_32, n_143);
  nor NOR2_g2181(n_30, n_122, n_32);
  nor NOR2_g2188(n_133, n_21, n_29);
  nor NOR2_g2175(n_28, n_42, n_143);
  nand NAND2_g2177(n_27, n_45, n_16);
  nor NOR2_g2179(n_39, in[4], n_32);
  xnor XNOR2_g2185(n_47, n_20, n_37);
  not NOT1_g2189(n_35, n_143);
  xnor XNOR2_g2190(n_119, n_38, in[0]);
  xnor XNOR2_g2191(n_32, n_25, in[6]);
  xnor XNOR2_g2192(n_143, n_25, in[5]);
  nor NOR2_g2195(n_24, n_122, n_23);
  nor NOR2_g2196(n_29, in[5], n_23);
  xnor XNOR2_g2187(n_45, n_25, n_15);
  nor NOR2_g2193(n_21, n_4, n_38);
  nor NOR2_g2194(n_20, n_122, n_42);
  not NOT1_g2197(n_23, n_38);
  xnor XNOR2_g2201(n_128, n_19, n_9);
  xnor XNOR2_g2199(n_38, n_37, in[6]);
  xnor XNOR2_g2198(n_25, in[3], n_8);
  xnor XNOR2_g2200(n_42, n_19, n_13);
  not NOT1_g2202(n_16, n_122);
  xnor XNOR2_g2207(n_15, in[1], in[0]);
  xnor XNOR2_g2208(n_13, in[1], in[7]);
  xnor XNOR2_g2210(n_11, in[0], in[7]);
  xnor XNOR2_g2204(n_9, in[1], in[5]);
  xnor XNOR2_g2209(n_8, in[2], in[7]);
  xnor XNOR2_g2203(n_7, in[3], in[5]);
  xnor XNOR2_g2211(n_19, in[2], in[6]);
  xnor XNOR2_g2205(n_37, in[1], in[4]);
  xnor XNOR2_g2206(n_122, in[7], in[5]);
  not NOT1_g2225(n_4, in[5]);
endmodule

